module top_module (
    input  wire in,
    output wire out
);
    assign out = in;
endmodule
