module top_module (
    output wire out
);
    assign out = 1'b0;
endmodule
